always @(posedge i_cpu_clk) begin
    if (i_rst) begin
    end else if (delaying) begin
    end else if (cycle_1_6502) begin
    end else if (cycle_2_6502) begin
        if (op_80_BRA) begin 
        end else if (~op_33_WTX) begin
            `PC <= inc_pc;
        end
    end else if (cycle_3_6502) begin
        if (am_ABS_a) begin
            if (op_JMP | op_JSR) begin
                `PC <= {reg_bram_doa_r, `ADDR0};
            end
        end else if (~am_IMM_m) begin
            if (am_PCR_r) begin
                if (op_BBR | op_BBS) begin
                end else begin
                    `PC <= `PC + {(reg_address[7] ? `ONES_8 : `ZERO_8), `ADDR0};
                end
            end else if (~op_33_WTX) begin
                `PC <= inc_pc;
            end
        end
    end else if (cycle_5_6502) begin
        if (op_BBR) begin
            if ((wire_data_byte_0 & reg_which) == 0) begin
                `PC <= `PC + {(wire_data_byte_0[7] ? `ONES_8 : `ZERO_8), wire_data_byte_0};
            end
        end else if (op_BBS) begin
            if ((wire_data_byte_0 & reg_which) != 0) begin
                `PC <= `PC + {(wire_data_byte_0[7] ? `ONES_8 : `ZERO_8), wire_data_byte_0};
            end
        end
    end else if (cycle_6_6502) begin
        if (am_AIIX_A_X | am_AIA_A) begin
            if (op_JMP) begin
                `PC <= {wire_data_byte_0, `IADDR0};
            end
        end
    end else if (cycle_1_65832) begin
    end
end
