always @(posedge i_clk) begin
    if (i_rst) begin
        ame_AIX_a_x <= 0;
    end else if (delaying) begin
    end else if (cycle_1_65832) begin
    end
end
