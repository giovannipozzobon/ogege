always @(posedge i_rst or posedge i_clk) begin
    if (i_rst) begin
        ame_IMM_m <= 0;
    end else if (cycle_1_65832) begin
    end
end
