always @(posedge i_rst or posedge i_clk) begin
    if (i_rst) begin
        op_STZ <= 0;
    end else if (delaying) begin
    end else if (cycle_1_6502) begin
        if (op_64_STZ | op_74_STZ | op_9C_STZ | op_9E_STZ) begin
            op_STZ <= 1;
        end
    end else if (cycle_4_6502) begin
        if (am_ABS_a) begin
            op_STZ <= 0;
        end
    end else if (cycle_1_65832) begin
    end
end
